module adder_TB();
	reg [31:0]Number1, Number2;
	reg reset, clk;
	wire [31:0]Result;
	
	IEEE_SP_FP_ADDER ia1(clk,reset,Number1,Number2,Result);
	
	always 
	#2 clk = ~clk;
	
	initial begin
	#2 clk=1;
    reset=1;
        
       #4 reset=0;
           
    Number1 = 32'b0100_0010_1100_0110_0000_0000_0000_0000;   //99
	Number2 = 32'b0100_0011_0011_0010_0000_0000_0000_0000;   //178   */

    #4;Number1 = 32'b0100_0010_1100_0010_0000_0000_0000_0000;   //97
	Number2 = 32'b1100_0010_1001_1110_0000_0000_0000_0000;   //-79

    #4;Number1 = 32'b1100_0010_0101_1100_0000_0000_0000_0000;   //-55
	Number2 = 32'b0100_0010_1001_0110_0000_0000_0000_0000;   //75 
    #4;Number1 = 32'b1100_0011_1000_1100_0000_0000_0000_0000;   //-280
	Number2 = 32'b1100_0010_1000_1010_0000_0000_0000_0000;   //-69 
    #4;Number1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;   //0
	Number2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;   //0 
    #4;Number1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;   //0
	Number2 = 32'b1100_0010_1110_0010_0000_0000_0000_0000;   //-113 
    #2;
        
    #200 $finish;
	end

	initial begin
		$dumpfile("adder_test.vcd");
		$dumpvars(0,tieee);
	end
endmodule